module decryption ( 
    input  wire        clk,
    input  wire        rst,
    input  wire        start,
    input  wire [63:0] key,
    input  wire [63:0] ciphertext,
    output reg  [63:0] decryptedtext,
    output reg         DECRYPT_DONE
); // inputs declaration


    // registers
    reg [31:0] temp, left, right;

    reg [31:0] p_array [0:17];
    reg [31:0] s_box0  [0:255];
    reg [31:0] s_box1  [0:255];
    reg [31:0] s_box2  [0:255];
    reg [31:0] s_box3  [0:255];

    reg [4:0] round;
    reg [3:0] state;
    reg       init;


    // local parameter
    localparam IDLE             = 4'd0,
               INIT             = 4'd1,
               DECRYPTION_LEFT  = 4'd2,
               DECRYPTION_RIGHT = 4'd3,
               DONE             = 4'd4,
               ENCRYPT_UNDO     = 4'd5,
               TRANSITION       = 4'd6,
               DECRYPT_LEFT     = 4'd7,
               DECRYPT_RIGHT    = 4'd8;


    // F-function of 4 sbox
    function [31:0] F;
        input [31:0] x;
        begin
            F = ( (s_box0[x[31:24]] + s_box1[x[23:16]]) ^
                  (s_box2[x[15:8]]) ) +
                  (s_box3[x[7:0]]);
        end
    endfunction


    // FSM logic
    always @(posedge clk) begin
        if (rst) begin

			//$readmemh("p_array.hex",p_array);
			//$readmemh("sbox0.hex",s_box0);
		  //$readmemh("sbox1.hex",s_box1);
			//$readmemh("sbox2.hex",s_box2);
			//$readmemh("sbox3.hex",s_box3);
		  
                  
			//insert p-array here
			p_array[0]  <= 32'h243f6a88;
			p_array[1]  <= 32'h85a308d3;
			p_array[2]  <= 32'h13198a2e;
			p_array[3]  <= 32'h03707344;
			p_array[4]  <= 32'ha4093822;
			p_array[5]  <= 32'h299f31d0;
			p_array[6]  <= 32'h082efa98;
			p_array[7]  <= 32'hec4e6c89;
			p_array[8]  <= 32'h452821e6;
			p_array[9]  <= 32'h38d01377;
			p_array[10] <= 32'hbe5466cf;
			p_array[11] <= 32'h34e90c6c;
			p_array[12] <= 32'hc0ac29b7;
			p_array[13] <= 32'hc97c50dd;
			p_array[14] <= 32'h3f84d5b5;
			p_array[15] <= 32'hb5470917;
			p_array[16] <= 32'h9216d5d9;
			p_array[17] <= 32'h8979fb1b;
			
			// sbox 0
			s_box0[0] <= 32'hd1310ba6;
			s_box0[1] <= 32'h98dfb5ac;
			s_box0[2] <= 32'h2ffd72db;
			s_box0[3] <= 32'hd01adfb7;
			s_box0[4] <= 32'hb8e1afed;
			s_box0[5] <= 32'h6a267e96;
			s_box0[6] <= 32'hba7c9045;
			s_box0[7] <= 32'hf12c7f99;
			s_box0[8] <= 32'h24a19947;
			s_box0[9] <= 32'hb3916cf7;
			s_box0[10] <= 32'h0801f2e2;
			s_box0[11] <= 32'h858efc16;
			s_box0[12] <= 32'h636920d8;
			s_box0[13] <= 32'h71574e69;
			s_box0[14] <= 32'ha458fea3;
			s_box0[15] <= 32'hf4933d7e;
			s_box0[16] <= 32'h0d95748f;
			s_box0[17] <= 32'h728eb658;
			s_box0[18] <= 32'h718bcd58;
			s_box0[19] <= 32'h82154aee;
			s_box0[20] <= 32'h7b54a41d;
			s_box0[21] <= 32'hc25a59b5;
			s_box0[22] <= 32'h9c30d539;
			s_box0[23] <= 32'h2af26013;
			s_box0[24] <= 32'hc5d1b023;
			s_box0[25] <= 32'h286085f0;
			s_box0[26] <= 32'hca417918;
			s_box0[27] <= 32'hb8db38ef;
			s_box0[28] <= 32'h8e79dcb0;
			s_box0[29] <= 32'h603a180e;
			s_box0[30] <= 32'h6c9e0e8b;
			s_box0[31] <= 32'hb01e8a3e;
			s_box0[32] <= 32'hd71577c1;
			s_box0[33] <= 32'hbd314b27;
			s_box0[34] <= 32'h78af2fda;
			s_box0[35] <= 32'h55605c60;
			s_box0[36] <= 32'he65525f3;
			s_box0[37] <= 32'haa55ab94;
			s_box0[38] <= 32'h57489862;
			s_box0[39] <= 32'h63e81440;
			s_box0[40] <= 32'h55ca396a;
			s_box0[41] <= 32'h2aab10b6;
			s_box0[42] <= 32'hb4cc5c34;
			s_box0[43] <= 32'h1141e8ce;
			s_box0[44] <= 32'ha15486af;
			s_box0[45] <= 32'h7c72e993;
			s_box0[46] <= 32'hb3ee1411;
			s_box0[47] <= 32'h636fbc2a;
			s_box0[48] <= 32'h2ba9c55d;
			s_box0[49] <= 32'h741831f6;
			s_box0[50] <= 32'hce5c3e16;
			s_box0[51] <= 32'h9b87931e;
			s_box0[52] <= 32'hafd6ba33;
			s_box0[53] <= 32'h6c24cf5c;
			s_box0[54] <= 32'h7a325381;
			s_box0[55] <= 32'h28958677;
			s_box0[56] <= 32'h3b8f4898;
			s_box0[57] <= 32'h6b4bb9af;
			s_box0[58] <= 32'hc4bfe81b;
			s_box0[59] <= 32'h66282193;
			s_box0[60] <= 32'h61d809cc;
			s_box0[61] <= 32'hfb21a991;
			s_box0[62] <= 32'h487cac60;
			s_box0[63] <= 32'h5dec8032;
			s_box0[64] <= 32'hef845d5d;
			s_box0[65] <= 32'he98575b1;
			s_box0[66] <= 32'hdc262302;
			s_box0[67] <= 32'heb651b88;
			s_box0[68] <= 32'h23893e81;
			s_box0[69] <= 32'hd396acc5;
			s_box0[70] <= 32'h0f6d6ff3;
			s_box0[71] <= 32'h83f44239;
			s_box0[72] <= 32'h2e0b4482;
			s_box0[73] <= 32'ha4842004;
			s_box0[74] <= 32'h69c8f04a;
			s_box0[75] <= 32'h9e1f9b5e;
			s_box0[76] <= 32'h21c66842;
			s_box0[77] <= 32'hf6e96c9a;
			s_box0[78] <= 32'h670c9c61;
			s_box0[79] <= 32'habd388f0;
			s_box0[80] <= 32'h6a51a0d2;
			s_box0[81] <= 32'hd8542f68;
			s_box0[82] <= 32'h960fa728;
			s_box0[83] <= 32'hab5133a3;
			s_box0[84] <= 32'h6eef0b6c;
			s_box0[85] <= 32'h137a3be4;
			s_box0[86] <= 32'hba3bf050;
			s_box0[87] <= 32'h7efb2a98;
			s_box0[88] <= 32'ha1f1651d;
			s_box0[89] <= 32'h39af0176;
			s_box0[90] <= 32'h66ca593e;
			s_box0[91] <= 32'h82430e88;
			s_box0[92] <= 32'h8cee8619;
			s_box0[93] <= 32'h456f9fb4;
			s_box0[94] <= 32'h7d84a5c3;
			s_box0[95] <= 32'h3b8b5ebe;
			s_box0[96] <= 32'he06f75d8;
			s_box0[97] <= 32'h85c12073;
			s_box0[98] <= 32'h401a449f;
			s_box0[99] <= 32'h56c16aa6;
			s_box0[100] <= 32'h4ed3aa62;
			s_box0[101] <= 32'h363f7706;
			s_box0[102] <= 32'h1bfedf72;
			s_box0[103] <= 32'h429b023d;
			s_box0[104] <= 32'h37d0d724;
			s_box0[105] <= 32'hd00a1248;
			s_box0[106] <= 32'hdb0fead3;
			s_box0[107] <= 32'h49f1c09b;
			s_box0[108] <= 32'h075372c9;
			s_box0[109] <= 32'h80991b7b;
			s_box0[110] <= 32'h25d479d8;
			s_box0[111] <= 32'hf6e8def7;
			s_box0[112] <= 32'he3fe501a;
			s_box0[113] <= 32'hb6794c3b;
			s_box0[114] <= 32'h976ce0bd;
			s_box0[115] <= 32'h04c006ba;
			s_box0[116] <= 32'hc1a94fb6;
			s_box0[117] <= 32'h409f60c4;
			s_box0[118] <= 32'h5e5c9ec2;
			s_box0[119] <= 32'h196a2463;
			s_box0[120] <= 32'h68fb6faf;
			s_box0[121] <= 32'h3e6c53b5;
			s_box0[122] <= 32'h1339b2eb;
			s_box0[123] <= 32'h3b52ec6f;
			s_box0[124] <= 32'h6dfc511f;
			s_box0[125] <= 32'h9b30952c;
			s_box0[126] <= 32'hcc814544;
			s_box0[127] <= 32'haf5ebd09;
			s_box0[128] <= 32'hbee3d004;
			s_box0[129] <= 32'hde334afd;
			s_box0[130] <= 32'h660f2807;
			s_box0[131] <= 32'h192e4bb3;
			s_box0[132] <= 32'hc0cba857;
			s_box0[133] <= 32'h45c8740f;
			s_box0[134] <= 32'hd20b5f39;
			s_box0[135] <= 32'hb9d3fbdb;
			s_box0[136] <= 32'h5579c0bd;
			s_box0[137] <= 32'h1a60320a;
			s_box0[138] <= 32'hd6a100c6;
			s_box0[139] <= 32'h402c7279;
			s_box0[140] <= 32'h679f25fe;
			s_box0[141] <= 32'hfb1fa3cc;
			s_box0[142] <= 32'h8ea5e9f8;
			s_box0[143] <= 32'hdb3222f8;
			s_box0[144] <= 32'h3c7516df;
			s_box0[145] <= 32'hfd616b15;
			s_box0[146] <= 32'h2f501ec8;
			s_box0[147] <= 32'had0552ab;
			s_box0[148] <= 32'h323db5fa;
			s_box0[149] <= 32'hfd238760;
			s_box0[150] <= 32'h53317b48;
			s_box0[151] <= 32'h3e00df82;
			s_box0[152] <= 32'h9e5c57bb;
			s_box0[153] <= 32'hca6f8ca0;
			s_box0[154] <= 32'h1a87562e;
			s_box0[155] <= 32'hdf1769db;
			s_box0[156] <= 32'hd542a8f6;
			s_box0[157] <= 32'h287effc3;
			s_box0[158] <= 32'hac6732c6;
			s_box0[159] <= 32'h8c4f5573;
			s_box0[160] <= 32'h695b27b0;
			s_box0[161] <= 32'hbbca58c8;
			s_box0[162] <= 32'he1ffa35d;
			s_box0[163] <= 32'hb8f011a0;
			s_box0[164] <= 32'h10fa3d98;
			s_box0[165] <= 32'hfd2183b8;
			s_box0[166] <= 32'h4afcb56c;
			s_box0[167] <= 32'h2dd1d35b;
			s_box0[168] <= 32'h9a53e479;
			s_box0[169] <= 32'hb6f84565;
			s_box0[170] <= 32'hd28e49bc;
			s_box0[171] <= 32'h4bfb9790;
			s_box0[172] <= 32'he1ddf2da;
			s_box0[173] <= 32'ha4cb7e33;
			s_box0[174] <= 32'h62fb1341;
			s_box0[175] <= 32'hcee4c6e8;
			s_box0[176] <= 32'hef20cada;
			s_box0[177] <= 32'h36774c01;
			s_box0[178] <= 32'hd07e9efe;
			s_box0[179] <= 32'h2bf11fb4;
			s_box0[180] <= 32'h95dbda4d;
			s_box0[181] <= 32'hae909198;
			s_box0[182] <= 32'heaad8e71;
			s_box0[183] <= 32'h6b93d5a0;
			s_box0[184] <= 32'hd08ed1d0;
			s_box0[185] <= 32'hafc725e0;
			s_box0[186] <= 32'h8e3c5b2f;
			s_box0[187] <= 32'h8e7594b7;
			s_box0[188] <= 32'h8ff6e2fb;
			s_box0[189] <= 32'hf2122b64;
			s_box0[190] <= 32'h8888b812;
			s_box0[191] <= 32'h900df01c;
			s_box0[192] <= 32'h4fad5ea0;
			s_box0[193] <= 32'h688fc31c;
			s_box0[194] <= 32'hd1cff191;
			s_box0[195] <= 32'hb3a8c1ad;
			s_box0[196] <= 32'h2f2f2218;
			s_box0[197] <= 32'hbe0e1777;
			s_box0[198] <= 32'hea752dfe;
			s_box0[199] <= 32'h8b021fa1;
			s_box0[200] <= 32'he5a0cc0f;
			s_box0[201] <= 32'hb56f74e8;
			s_box0[202] <= 32'h18acf3d6;
			s_box0[203] <= 32'hce89e299;
			s_box0[204] <= 32'hb4a84fe0;
			s_box0[205] <= 32'hfd13e0b7;
			s_box0[206] <= 32'h7cc43b81;
			s_box0[207] <= 32'hd2ada8d9;
			s_box0[208] <= 32'h165fa266;
			s_box0[209] <= 32'h80957705;
			s_box0[210] <= 32'h93cc7314;
			s_box0[211] <= 32'h211a1477;
			s_box0[212] <= 32'he6ad2065;
			s_box0[213] <= 32'h77b5fa86;
			s_box0[214] <= 32'hc75442f5;
			s_box0[215] <= 32'hfb9d35cf;
			s_box0[216] <= 32'hebcdaf0c;
			s_box0[217] <= 32'h7b3e89a0;
			s_box0[218] <= 32'hd6411bd3;
			s_box0[219] <= 32'hae1e7e49;
			s_box0[220] <= 32'h00250e2d;
			s_box0[221] <= 32'h2071b35e;
			s_box0[222] <= 32'h226800bb;
			s_box0[223] <= 32'h57b8e0af;
			s_box0[224] <= 32'h2464369b;
			s_box0[225] <= 32'hf009b91e;
			s_box0[226] <= 32'h5563911d;
			s_box0[227] <= 32'h59dfa6aa;
			s_box0[228] <= 32'h78c14389;
			s_box0[229] <= 32'hd95a537f;
			s_box0[230] <= 32'h207d5ba2;
			s_box0[231] <= 32'h02e5b9c5;
			s_box0[232] <= 32'h83260376;
			s_box0[233] <= 32'h6295cfa9;
			s_box0[234] <= 32'h11c81968;
			s_box0[235] <= 32'h4e734a41;
			s_box0[236] <= 32'hb3472dca;
			s_box0[237] <= 32'h7b14a94a;
			s_box0[238] <= 32'h1b510052;
			s_box0[239] <= 32'h9a532915;
			s_box0[240] <= 32'hd60f573f;
			s_box0[241] <= 32'hbc9bc6e4;
			s_box0[242] <= 32'h2b60a476;
			s_box0[243] <= 32'h81e67400;
			s_box0[244] <= 32'h08ba6fb5;
			s_box0[245] <= 32'h571be91f;
			s_box0[246] <= 32'hf296ec6b;
			s_box0[247] <= 32'h2a0dd915;
			s_box0[248] <= 32'hb6636521;
			s_box0[249] <= 32'he7b9f9b6;
			s_box0[250] <= 32'hff34052e;
			s_box0[251] <= 32'hc5855664;
			s_box0[252] <= 32'h53b02d5d;
			s_box0[253] <= 32'ha99f8fa1;
			s_box0[254] <= 32'h08ba4799;
			s_box0[255] <= 32'h6e85076a;
			
			// sbox 1			problem
			s_box1[0]   <= 32'h4b7a70e9;
			s_box1[1]   <= 32'hb5b32944;
			s_box1[2]   <= 32'hdb75092e;
			s_box1[3]   <= 32'hc4192623;
			s_box1[4]   <= 32'had6ea6b0;
			s_box1[5]   <= 32'h49a7df7d;
			s_box1[6]   <= 32'h9cee60b8;
			s_box1[7]   <= 32'h8fedb266;
			s_box1[8]   <= 32'hecaa8c71;
			s_box1[9]   <= 32'h699a17ff;
			s_box1[10]  <= 32'h5664526c;
			s_box1[11]  <= 32'hc2b19ee1;
			s_box1[12]  <= 32'h193602a5;
			s_box1[13]  <= 32'h75094c29;
			s_box1[14]  <= 32'ha0591340;
			s_box1[15]  <= 32'he4183a3e;
			s_box1[16]  <= 32'h3f54989a;
			s_box1[17]  <= 32'h5b429d65;
			s_box1[18]  <= 32'h6b8fe4d6;
			s_box1[19]  <= 32'h99f73fd6;
			s_box1[20]  <= 32'ha1d29c07;
			s_box1[21]  <= 32'hefe830f5;
			s_box1[22]  <= 32'h4d2d38e6;
			s_box1[23]  <= 32'hf0255dc1;
			s_box1[24]  <= 32'h4cdd2086;
			s_box1[25]  <= 32'h8470eb26;
			s_box1[26]  <= 32'h6382e9c6;
			s_box1[27]  <= 32'h021ecc5e;
			s_box1[28]  <= 32'h09686b3f;
			s_box1[29]  <= 32'h3ebaefc9;
			s_box1[30]  <= 32'h3c971814;
			s_box1[31]  <= 32'h6b6a70a1;
			s_box1[32]  <= 32'h687f3584;
			s_box1[33]  <= 32'h52a0e286;
			s_box1[34]  <= 32'hb79c5305;
			s_box1[35]  <= 32'haa500737;
			s_box1[36]  <= 32'h3e07841c;
			s_box1[37]  <= 32'h7fdeae5c;
			s_box1[38]  <= 32'h8e7d44ec;
			s_box1[39]  <= 32'h5716f2b8;
			s_box1[40]  <= 32'hb03ada37;
			s_box1[41]  <= 32'hf0500c0d;
			s_box1[42]  <= 32'hf01c1f04;
			s_box1[43]  <= 32'h0200b3ff;
			s_box1[44]  <= 32'hae0cf51a;
			s_box1[45]  <= 32'h3cb574b2;
			s_box1[46]  <= 32'h25837a58;
			s_box1[47]  <= 32'hdc0921bd;
			s_box1[48]  <= 32'hd19113f9;
			s_box1[49]  <= 32'h7ca92ff6;
			s_box1[50]  <= 32'h94324773;
			s_box1[51]  <= 32'h22f54701;
			s_box1[52]  <= 32'h3ae5e581;
			s_box1[53]  <= 32'h37c2dadc;
			s_box1[54]  <= 32'hc8b57634;
			s_box1[55]  <= 32'h9af3dda7;
			s_box1[56]  <= 32'ha9446146;
			s_box1[57]  <= 32'h0fd0030e;
			s_box1[58]  <= 32'hecc8c73e;
			s_box1[59]  <= 32'ha4751e41;
			s_box1[60]  <= 32'he238cd99;
			s_box1[61]  <= 32'h3bea0e2f;
			s_box1[62]  <= 32'h3280bba1;
			s_box1[63]  <= 32'h183eb331;
			s_box1[64]  <= 32'h4e548b38;
			s_box1[65]  <= 32'h4f6db908;
			s_box1[66]  <= 32'h6f420d03;
			s_box1[67]  <= 32'hf60a04bf;
			s_box1[68]  <= 32'h2cb81290;
			s_box1[69]  <= 32'h24977c79;
			s_box1[70]  <= 32'h5679b072;
			s_box1[71]  <= 32'hbcaf89af;
			s_box1[72]  <= 32'hde9a771f;
			s_box1[73]  <= 32'hd9930810;
			s_box1[74]  <= 32'hb38bae12;
			s_box1[75]  <= 32'hdccf3f2e;
			s_box1[76]  <= 32'h5512721f;
			s_box1[77]  <= 32'h2e6b7124;
			s_box1[78]  <= 32'h501adde6;
			s_box1[79]  <= 32'h9f84cd87;
			s_box1[80]  <= 32'h7a584718;
			s_box1[81]  <= 32'h7408da17;
			s_box1[82]  <= 32'hbc9f9abc;
			s_box1[83]  <= 32'he94b7d8c;
			s_box1[84]  <= 32'hec7aec3a;
			s_box1[85]  <= 32'hdb851dfa;
			s_box1[86]  <= 32'h63094366;
			s_box1[87]  <= 32'hc464c3d2;
			s_box1[88]  <= 32'hef1c1847;
			s_box1[89]  <= 32'h3215d908;
			s_box1[90]  <= 32'hdd433b37;
			s_box1[91]  <= 32'h24c2ba16;
			s_box1[92]  <= 32'h12a14d43;
			s_box1[93]  <= 32'h2a65c451;
			s_box1[94]  <= 32'h50940002;
			s_box1[95]  <= 32'h133ae4dd;
			s_box1[96]  <= 32'h71dff89e;
			s_box1[97]  <= 32'h10314e55;
			s_box1[98]  <= 32'h81ac77d6;
			s_box1[99]  <= 32'h5f11199b;
			s_box1[100] <= 32'h043556f1;
			s_box1[101] <= 32'hd7a3c76b;
			s_box1[102] <= 32'h3c11183b;
			s_box1[103] <= 32'h5924a509;
			s_box1[104] <= 32'hf28fe6ed;
			s_box1[105] <= 32'h97f1fbfa;
			s_box1[106] <= 32'h9ebabf2c;
			s_box1[107] <= 32'h1e153c6e;
			s_box1[108] <= 32'h86e34570;
			s_box1[109] <= 32'heae96fb1;
			s_box1[110] <= 32'h860e5e0a;
			s_box1[111] <= 32'h5a3e2ab3;
			s_box1[112] <= 32'h771fe71c;
			s_box1[113] <= 32'h4e3d06fa;
			s_box1[114] <= 32'h2965dcb9;
			s_box1[115] <= 32'h99e71d0f;
			s_box1[116] <= 32'h803e89d6;
			s_box1[117] <= 32'h5266c825;
			s_box1[118] <= 32'h2e4cc978;
			s_box1[119] <= 32'h9c10b36a;
			s_box1[120] <= 32'hc6150eba;
			s_box1[121] <= 32'h94e2ea78;
			s_box1[122] <= 32'ha5fc3c53;
			s_box1[123] <= 32'h1e0a2df4;
			s_box1[124] <= 32'hf2f74ea7;
			s_box1[125] <= 32'h361d2b3d;
			s_box1[126] <= 32'h1939260f;
			s_box1[127] <= 32'h19c27960;
			s_box1[128] <= 32'h5223a708;
			s_box1[129] <= 32'hf71312b6;
			s_box1[130] <= 32'hebadfe6e;
			s_box1[131] <= 32'heac31f66;
			s_box1[132] <= 32'he3bc4595;
			s_box1[133] <= 32'ha67bc883;
			s_box1[134] <= 32'hb17f37d1;
			s_box1[135] <= 32'h018cff28;
			s_box1[136] <= 32'hc332ddef;
			s_box1[137] <= 32'hbe6c5aa5;
			s_box1[138] <= 32'h65582185;
			s_box1[139] <= 32'h68ab9802;
			s_box1[140] <= 32'heecea50f;
			s_box1[141] <= 32'hdb2f953b;
			s_box1[142] <= 32'h2aef7dad;
			s_box1[143] <= 32'h5b6e2f84;
			s_box1[144] <= 32'h1521b628;
			s_box1[145] <= 32'h29076170;
			s_box1[146] <= 32'hecdd4775;
			s_box1[147] <= 32'h619f1510;
			s_box1[148] <= 32'h13cca830;
			s_box1[149] <= 32'heb61bd96;
			s_box1[150] <= 32'h0334fe1e;
			s_box1[151] <= 32'haa0363cf;
			s_box1[152] <= 32'hb5735c90;
			s_box1[153] <= 32'h4c70a239;
			s_box1[154] <= 32'hd59e9e0b;
			s_box1[155] <= 32'hcbaade14;
			s_box1[156] <= 32'heecc86bc;
			s_box1[157] <= 32'h60622ca7;
			s_box1[158] <= 32'h9cab5cab;
			s_box1[159] <= 32'hb2f3846e;
			s_box1[160] <= 32'h648b1eaf;
			s_box1[161] <= 32'h19bdf0ca;
			s_box1[162] <= 32'ha02369b9;
			s_box1[163] <= 32'h655abb50;
			s_box1[164] <= 32'h40685a32;
			s_box1[165] <= 32'h3c2ab4b3;
			s_box1[166] <= 32'h319ee9d5;
			s_box1[167] <= 32'hc021b8f7;
			s_box1[168] <= 32'h9b540b19;
			s_box1[169] <= 32'h875fa099;
			s_box1[170] <= 32'h95f7997e;
			s_box1[171] <= 32'h623d7da8;
			s_box1[172] <= 32'hf837889a;
			s_box1[173] <= 32'h97e32d77;
			s_box1[174] <= 32'h11ed935f;
			s_box1[175] <= 32'h16681281;
			s_box1[176] <= 32'h0e358829;
			s_box1[177] <= 32'hc7e61fd6;
			s_box1[178] <= 32'h96dedfa1;
			s_box1[179] <= 32'h7858ba99;
			s_box1[180] <= 32'h57f584a5;
			s_box1[181] <= 32'h1b227263;
			s_box1[182] <= 32'h9b83c3ff;
			s_box1[183] <= 32'h1ac246e6;
			s_box1[184] <= 32'h7472dd37;
			s_box1[185] <= 32'h99451121;
			s_box1[186] <= 32'h91d90c91;
			s_box1[187] <= 32'h19069695;
			s_box1[188] <= 32'h40f98402;
			s_box1[189] <= 32'h7c14a84d;
			s_box1[190] <= 32'h3c49e798;
			s_box1[191] <= 32'h566538c7;
			s_box1[192] <= 32'h26868593;
			s_box1[193] <= 32'h98c08126;
			s_box1[194] <= 32'h2a36c92b;
			s_box1[195] <= 32'h68494101;
			s_box1[196] <= 32'h47652259;
			s_box1[197] <= 32'h8606f0e2;
			s_box1[198] <= 32'h5343b67e;
			s_box1[199] <= 32'h85a75892;
			s_box1[200] <= 32'h5f74f74d;
			s_box1[201] <= 32'h217c2a71;
			s_box1[202] <= 32'h706b4765;
			s_box1[203] <= 32'h321876e5;
			s_box1[204] <= 32'h96e7365c;
			s_box1[205] <= 32'h96b52815;
			s_box1[206] <= 32'h02919d67;
			s_box1[207] <= 32'h6f62b721;
			s_box1[208] <= 32'h322f9862;
			s_box1[209] <= 32'h9407760d;
			s_box1[210] <= 32'h875f12a2;
			s_box1[211] <= 32'h9674994d;
			s_box1[212] <= 32'h27f311c1;
			s_box1[213] <= 32'h445171af;
			s_box1[214]   <= 32'h0d09222c;
			s_box1[215]   <= 32'h986427b3;
			s_box1[216]   <= 32'h68962b8c;
			s_box1[217]   <= 32'h9f168f51;
			s_box1[218]   <= 32'h8ba8122c;
			s_box1[219]   <= 32'h15f33668;
			s_box1[220]   <= 32'h6109439f;
			s_box1[221]   <= 32'h991c4c16;
			s_box1[222]   <= 32'h07d9f783;
			s_box1[223]   <= 32'h9c762744;
			s_box1[224]  <= 32'h79949d1c;
			s_box1[225]  <= 32'h017596a7;
			s_box1[226]  <= 32'h74c803d9;
			s_box1[227]  <= 32'h2565615f;
			s_box1[228]  <= 32'h1d670606;
			s_box1[229]  <= 32'h69655928;
			s_box1[230]  <= 32'h70a8276f;
			s_box1[231]  <= 32'h5c246f91;
			s_box1[232]  <= 32'h5f69a528;
			s_box1[233]  <= 32'h8674995b;
			s_box1[234]  <= 32'h80d5d71c;
			s_box1[235]  <= 32'h5c197992;
			s_box1[236]  <= 32'h567922d3;
			s_box1[237]  <= 32'h5c3327d1;
			s_box1[238]  <= 32'h40c952c7;
			s_box1[239]  <= 32'h52a67744;
			s_box1[240]  <= 32'h6a908906;
			s_box1[241]  <= 32'h42636952;
			s_box1[242]  <= 32'h508a65b7;
			s_box1[243]  <= 32'h2499d7a2;
			s_box1[244]  <= 32'h7d922572;
			s_box1[245]  <= 32'h0491953f;
			s_box1[246]  <= 32'h52495c61;
			s_box1[247]  <= 32'h40c88599;
			s_box1[248]  <= 32'h7207aef0;
			s_box1[249]  <= 32'h98d169d5;
			s_box1[250]  <= 32'h45455a73;
			s_box1[251]  <= 32'h9658257a;
			s_box1[252]  <= 32'h089c8915;
			s_box1[253]  <= 32'h4223b24f;
			s_box1[254]  <= 32'h98c7e39a;
			s_box1[255]  <= 32'h2b96312a;

			//sbox 2
			s_box2[0] <= 32'h69002b28;
			s_box2[1] <= 32'h0764c2a5;
			s_box2[2] <= 32'h9980d8ef;
			s_box2[3] <= 32'hb5606c46;
			s_box2[4] <= 32'h6a47f017;
			s_box2[5] <= 32'h748f8241;
			s_box2[6] <= 32'h3c405621;
			s_box2[7] <= 32'h1c19b728;
			s_box2[8] <= 32'h4449830b;
			s_box2[9] <= 32'h74136eb1;
			s_box2[10] <= 32'h56d3969a;
			s_box2[11] <= 32'h04c97974;
			s_box2[12] <= 32'h1c7c25e2;
			s_box2[13] <= 32'h9661c5c3;
			s_box2[14] <= 32'h84118429;
			s_box2[15] <= 32'h15744b91;
			s_box2[16] <= 32'h6361c470;
			s_box2[17] <= 32'h9953c829;
			s_box2[18] <= 32'h7164995c;
			s_box2[19] <= 32'h6f68e92d;
			s_box2[20] <= 32'h4f91e921;
			s_box2[21] <= 32'h939622c5;
			s_box2[22] <= 32'h2f781912;
			s_box2[23] <= 32'h95b79607;
			s_box2[24] <= 32'h4634f591;
			s_box2[25] <= 32'h2f802183;
			s_box2[26] <= 32'h47738378;
			s_box2[27] <= 32'h669c5225;
			s_box2[28] <= 32'h2786960b;
			s_box2[29] <= 32'h715a3696;
			s_box2[30] <= 32'h65e31751;
			s_box2[31] <= 32'h82834b5b;
			s_box2[32] <= 32'h5721c0fc;
			s_box2[33] <= 32'h76162380;
			s_box2[34] <= 32'h4721a938;
			s_box2[35] <= 32'h42206c8b;
			s_box2[36] <= 32'h16f06762;
			s_box2[37] <= 32'h68925501;
			s_box2[38] <= 32'h4294025a;
			s_box2[39] <= 32'h44682dff;
			s_box2[40] <= 32'h7c87c073;
			s_box2[41] <= 32'h49c8642b;
			s_box2[42] <= 32'h8055938d;
			s_box2[43] <= 32'h534b0788;
			s_box2[44] <= 32'h2646f888;
			s_box2[45] <= 32'h97d8b589;
			s_box2[46] <= 32'h0623a65e;
			s_box2[47] <= 32'h79929117;
			s_box2[48] <= 32'h43e4811a;
			s_box2[49] <= 32'h82728952;
			s_box2[50] <= 32'h6479706b;
			s_box2[51] <= 32'h5164ab0c;
			s_box2[52] <= 32'h3c491102;
			s_box2[53] <= 32'h807095b9;
			s_box2[54] <= 32'h56860352;
			s_box2[55] <= 32'h61578f5a;
			s_box2[56] <= 32'h089c836c;
			s_box2[57] <= 32'h4f923c72;
			s_box2[58] <= 32'h4f989c1c;
			s_box2[59] <= 32'h5c6b4594;
			s_box2[60] <= 32'h27f29910;
			s_box2[61] <= 32'h21571217;
			s_box2[62] <= 32'h45455a73;
			s_box2[63] <= 32'h804d9561;
			s_box2[64] <= 32'h515792c8;
			s_box2[65] <= 32'h567922d3;
			s_box2[66] <= 32'h706b4765;
			s_box2[67] <= 32'h5a2971d5;
			s_box2[68] <= 32'h5f74f74d;
			s_box2[69] <= 32'h82728952;
			s_box2[70] <= 32'h217c2a71;
			s_box2[71] <= 32'h321876e5;
			s_box2[72] <= 32'h96e7365c;
			s_box2[73] <= 32'h96b52815;
			s_box2[74] <= 32'h02919d67;
			s_box2[75] <= 32'h6f62b721;
			s_box2[76] <= 32'h322f9862;
			s_box2[77] <= 32'h9407760d;
			s_box2[78] <= 32'h875f12a2;
			s_box2[79] <= 32'h9674994d;
			s_box2[80] <= 32'h27f311c1;
			s_box2[81] <= 32'h445171af;
			s_box2[82] <= 32'h0d09222c;
			s_box2[83] <= 32'h986427b3;
			s_box2[84] <= 32'h68962b8c;
			s_box2[85] <= 32'h9f168f51;
			s_box2[86] <= 32'h8ba8122c;
			s_box2[87] <= 32'h15f33668;
			s_box2[88] <= 32'h6109439f;
			s_box2[89] <= 32'h991c4c16;
			s_box2[90] <= 32'h07d9f783;
			s_box2[91] <= 32'h9c762744;
			s_box2[92] <= 32'h79949d1c;
			s_box2[93] <= 32'h017596a7;
			s_box2[94] <= 32'h74c803d9;
			s_box2[95] <= 32'h2565615f;
			s_box2[96] <= 32'h1d670606;
			s_box2[97] <= 32'h69655928;
			s_box2[98] <= 32'h70a8276f;
			s_box2[99] <= 32'h5c246f91;
			s_box2[100] <= 32'h5f69a528;
			s_box2[101] <= 32'h8674995b;
			s_box2[102] <= 32'h80d5d71c;
			s_box2[103] <= 32'h5c197992;
			s_box2[104] <= 32'h567922d3;
			s_box2[105] <= 32'h5c3327d1;
			s_box2[106] <= 32'h40c952c7;
			s_box2[107] <= 32'h52a67744;
			s_box2[108] <= 32'h6a908906;
			s_box2[109] <= 32'h42636952;
			s_box2[110] <= 32'h508a65b7;
			s_box2[111] <= 32'h2499d7a2;
			s_box2[112] <= 32'h7d922572;
			s_box2[113] <= 32'h0491953f;
			s_box2[114] <= 32'h52495c61;
			s_box2[115] <= 32'h40c88599;
			s_box2[116] <= 32'h7207aef0;
			s_box2[117] <= 32'h98d169d5;
			s_box2[118] <= 32'h45455a73;
			s_box2[119] <= 32'h9658257a;
			s_box2[120] <= 32'h089c8915;
			s_box2[121] <= 32'h4223b24f;
			s_box2[122] <= 32'h98c7e39a;
			s_box2[123] <= 32'h2b96312a;
			s_box2[124] <= 32'h69002b28;
			s_box2[125] <= 32'h0764c2a5;
			s_box2[126] <= 32'h9980d8ef;
			s_box2[127] <= 32'hb5606c46;
			s_box2[128] <= 32'h6a47f017;
			s_box2[129] <= 32'h748f8241;
			s_box2[130] <= 32'h3c405621;
			s_box2[131] <= 32'h1c19b728;
			s_box2[132] <= 32'h4449830b;
			s_box2[133] <= 32'h74136eb1;
			s_box2[134] <= 32'h56d3969a;
			s_box2[135] <= 32'h04c97974;
			s_box2[136] <= 32'h1c7c25e2;
			s_box2[137] <= 32'h9661c5c3;
			s_box2[138] <= 32'h84118429;
			s_box2[139] <= 32'h15744b91;
			s_box2[140] <= 32'h6361c470;
			s_box2[141] <= 32'h9953c829;
			s_box2[142] <= 32'h7164995c;
			s_box2[143] <= 32'h6f68e92d;
			s_box2[144] <= 32'h4f91e921;
			s_box2[145] <= 32'h939622c5;
			s_box2[146] <= 32'h2f781912;
			s_box2[147] <= 32'h95b79607;
			s_box2[148] <= 32'h4634f591;
			s_box2[149] <= 32'h2f802183;
			s_box2[150] <= 32'h47738378;
			s_box2[151] <= 32'h669c5225;
			s_box2[152] <= 32'h2786960b;
			s_box2[153] <= 32'h715a3696;
			s_box2[154] <= 32'h65e31751;
			s_box2[155] <= 32'h82834b5b;
			s_box2[156] <= 32'h5721c0fc;
			s_box2[157] <= 32'h76162380;
			s_box2[158] <= 32'h4721a938;
			s_box2[159] <= 32'h42206c8b;
			s_box2[160] <= 32'h16f06762;
			s_box2[161] <= 32'h68925501;
			s_box2[162] <= 32'h4294025a;
			s_box2[163] <= 32'h44682dff;
			s_box2[164] <= 32'h7c87c073;
			s_box2[165] <= 32'h49c8642b;
			s_box2[166] <= 32'h8055938d;
			s_box2[167] <= 32'h534b0788;
			s_box2[168] <= 32'h2646f888;
			s_box2[169] <= 32'h97d8b589;
			s_box2[170] <= 32'h0623a65e;
			s_box2[171] <= 32'h79929117;
			s_box2[172] <= 32'h43e4811a;
			s_box2[173] <= 32'h82728952;
			s_box2[174] <= 32'h6479706b;
			s_box2[175] <= 32'h5164ab0c;
			s_box2[176] <= 32'h3c491102;
			s_box2[177] <= 32'h807095b9;
			s_box2[178] <= 32'h56860352;
			s_box2[179] <= 32'h61578f5a;
			s_box2[180] <= 32'h089c836c;
			s_box2[181] <= 32'h4f923c72;
			s_box2[182] <= 32'h4f989c1c;
			s_box2[183] <= 32'h5c6b4594;
			s_box2[184] <= 32'h27f29910;
			s_box2[185] <= 32'h21571217;
			s_box2[186] <= 32'h45455a73;
			s_box2[187] <= 32'h804d9561;
			s_box2[188] <= 32'h515792c8;
			s_box2[189] <= 32'h567922d3;
			s_box2[190] <= 32'h706b4765;
			s_box2[191] <= 32'h5a2971d5;
			s_box2[192] <= 32'h5f74f74d;
			s_box2[193] <= 32'h82728952;
			s_box2[194] <= 32'h217c2a71;
			s_box2[195] <= 32'h321876e5;
			s_box2[196] <= 32'h96e7365c;
			s_box2[197] <= 32'h96b52815;
			s_box2[198] <= 32'h02919d67;
			s_box2[199] <= 32'h6f62b721;
			s_box2[200] <= 32'h322f9862;
			s_box2[201] <= 32'h9407760d;
			s_box2[202] <= 32'h875f12a2;
			s_box2[203] <= 32'h9674994d;
			s_box2[204] <= 32'h27f311c1;
			s_box2[205] <= 32'h445171af;
			s_box2[206] <= 32'h0d09222c;
			s_box2[207] <= 32'h986427b3;
			s_box2[208] <= 32'h68962b8c;
			s_box2[209] <= 32'h9f168f51;
			s_box2[210] <= 32'h8ba8122c;
			s_box2[211] <= 32'h15f33668;
			s_box2[212] <= 32'h6109439f;
			s_box2[213] <= 32'h991c4c16;
			s_box2[214] <= 32'h07d9f783;
			s_box2[215] <= 32'h9c762744;
			s_box2[216] <= 32'h79949d1c;
			s_box2[217] <= 32'h017596a7;
			s_box2[218] <= 32'h74c803d9;
			s_box2[219] <= 32'h2565615f;
			s_box2[220] <= 32'h1d670606;
			s_box2[221] <= 32'h69655928;
			s_box2[222] <= 32'h70a8276f;
			s_box2[223] <= 32'h5c246f91;
			s_box2[224] <= 32'h5f69a528;
			s_box2[225] <= 32'h8674995b;
			s_box2[226] <= 32'h80d5d71c;
			s_box2[227] <= 32'h5c197992;
			s_box2[228] <= 32'h567922d3;
			s_box2[229] <= 32'h5c3327d1;
			s_box2[230] <= 32'h40c952c7;
			s_box2[231] <= 32'h52a67744;
			s_box2[232] <= 32'h6a908906;
			s_box2[233] <= 32'h42636952;
			s_box2[234] <= 32'h508a65b7;
			s_box2[235] <= 32'h2499d7a2;
			s_box2[236] <= 32'h7d922572;
			s_box2[237] <= 32'h0491953f;
			s_box2[238] <= 32'h52495c61;
			s_box2[239] <= 32'h40c88599;
			s_box2[240] <= 32'h7207aef0;
			s_box2[241] <= 32'h98d169d5;
			s_box2[242] <= 32'h45455a73;
			s_box2[243] <= 32'h9658257a;
			s_box2[244] <= 32'h089c8915;
			s_box2[245] <= 32'h4223b24f;
			s_box2[246] <= 32'h98c7e39a;
			s_box2[247] <= 32'h2b96312a;
			s_box2[248] <= 32'h69002b28;
			s_box2[249] <= 32'h0764c2a5;
			s_box2[250] <= 32'h9980d8ef;
			s_box2[251] <= 32'hb5606c46;
			s_box2[252] <= 32'h6a47f017;
			s_box2[253] <= 32'h748f8241;
			s_box2[254] <= 32'h3c405621;
			s_box2[255] <= 32'h1c19b728;
			
			//sbox 3
			s_box3[0]<= 32'h75b63e79;
			s_box3[1]<= 32'h58bfb5a0;
			s_box3[2]<= 32'h9750c3a9;
			s_box3[3]<= 32'h22c8c459;
			s_box3[4]<= 32'h76b32549;
			s_box3[5]<= 32'h8cdc3a36;
			s_box3[6]<= 32'h89151608;
			s_box3[7]<= 32'h2f87c582;
			s_box3[8]<= 32'h196291b1;
			s_box3[9]<= 32'h5b056ef8;
			s_box3[10]<= 32'h9c7a08b5;
			s_box3[11]<= 32'h84c8515f;
			s_box3[12]<= 32'h0d62b95b;
			s_box3[13]<= 32'h662a0c71;
			s_box3[14]<= 32'h56722237;
			s_box3[15]<= 32'h6f5f849c;
			s_box3[16]<= 32'h262a3641;
			s_box3[17]<= 32'h4b34b631;
			s_box3[18]<= 32'h4f923c72;
			s_box3[19]<= 32'h4f989c1c;
			s_box3[20]<= 32'h5c6b4594;
			s_box3[21]<= 32'h27f29910;
			s_box3[22]<= 32'h21571217;
			s_box3[23]<= 32'h45455a73;
			s_box3[24]<= 32'h804d9561;
			s_box3[25]<= 32'h515792c8;
			s_box3[26]<= 32'h567922d3;
			s_box3[27]<= 32'h706b4765;
			s_box3[28]<= 32'h5a2971d5;
			s_box3[29]<= 32'h5f74f74d;
			s_box3[30]<= 32'h82728952;
			s_box3[31]<= 32'h217c2a71;
			s_box3[32]<= 32'h321876e5;
			s_box3[33]<= 32'h96e7365c;
			s_box3[34]<= 32'h96b52815;
			s_box3[35]<= 32'h02919d67;
			s_box3[36]<= 32'h6f62b721;
			s_box3[37]<= 32'h322f9862;
			s_box3[38]<= 32'h9407760d;
			s_box3[39]<= 32'h875f12a2;
			s_box3[40]<= 32'h9674994d;
			s_box3[41]<= 32'h27f311c1;
			s_box3[42]<= 32'h445171af;
			s_box3[43]<= 32'h0d09222c;
			s_box3[44]<= 32'h986427b3;
			s_box3[45]<= 32'h68962b8c;
			s_box3[46]<= 32'h9f168f51;
			s_box3[47]<= 32'h8ba8122c;
			s_box3[48]<= 32'h15f33668;
			s_box3[49]<= 32'h6109439f;
			s_box3[50]<= 32'h991c4c16;
			s_box3[51]<= 32'h07d9f783;
			s_box3[52]<= 32'h9c762744;
			s_box3[53]<= 32'h79949d1c;
			s_box3[54]<= 32'h017596a7;
			s_box3[55]<= 32'h74c803d9;
			s_box3[56]<= 32'h2565615f;
			s_box3[57]<= 32'h1d670606;
			s_box3[58]<= 32'h69655928;
			s_box3[59]<= 32'h70a8276f;
			s_box3[60]<= 32'h5c246f91;
			s_box3[61]<= 32'h5f69a528;
			s_box3[62]<= 32'h8674995b;
			s_box3[63]<= 32'h80d5d71c;
			s_box3[64]<= 32'h5c197992;
			s_box3[65]<= 32'h567922d3;
			s_box3[66]<= 32'h5c3327d1;
			s_box3[67]<= 32'h40c952c7;
			s_box3[68]<= 32'h52a67744;
			s_box3[69]<= 32'h6a908906;
			s_box3[70]<= 32'h42636952;
			s_box3[71]<= 32'h508a65b7;
			s_box3[72]<= 32'h2499d7a2;
			s_box3[73]<= 32'h7d922572;
			s_box3[74]<= 32'h0491953f;
			s_box3[75]<= 32'h52495c61;
			s_box3[76]<= 32'h40c88599;
			s_box3[77]<= 32'h7207aef0;
			s_box3[78]<= 32'h98d169d5;
			s_box3[79]<= 32'h45455a73;
			s_box3[80]<= 32'h9658257a;
			s_box3[81]<= 32'h089c8915;
			s_box3[82]<= 32'h4223b24f;
			s_box3[83]<= 32'h98c7e39a;
			s_box3[84]<= 32'h2b96312a;
			s_box3[85]<= 32'h75b63e79;
			s_box3[86]<= 32'h58bfb5a0;
			s_box3[87]<= 32'h9750c3a9;
			s_box3[88]<= 32'h22c8c459;
			s_box3[89]<= 32'h76b32549;
			s_box3[90]<= 32'h8cdc3a36;
			s_box3[91]<= 32'h89151608;
			s_box3[92]<= 32'h2f87c582;
			s_box3[93]<= 32'h196291b1;
			s_box3[94]<= 32'h5b056ef8;
			s_box3[95]<= 32'h9c7a08b5;
			s_box3[96]<= 32'h84c8515f;
			s_box3[97]<= 32'h0d62b95b;
			s_box3[98]<= 32'h662a0c71;
			s_box3[99]<= 32'h56722237;
			s_box3[100]<= 32'h6f5f849c;
			s_box3[101]<= 32'h262a3641;
			s_box3[102]<= 32'h4b34b631;
			s_box3[103]<= 32'h4f923c72;
			s_box3[104]<= 32'h4f989c1c;
			s_box3[105]<= 32'h5c6b4594;
			s_box3[106]<= 32'h27f29910;
			s_box3[107]<= 32'h21571217;
			s_box3[108]<= 32'h45455a73;
			s_box3[109]<= 32'h804d9561;
			s_box3[110]<= 32'h515792c8;
			s_box3[111]<= 32'h567922d3;
			s_box3[112]<= 32'h706b4765;
			s_box3[113]<= 32'h5a2971d5;
			s_box3[114]<= 32'h5f74f74d;
			s_box3[115]<= 32'h82728952;
			s_box3[116]<= 32'h217c2a71;
			s_box3[117]<= 32'h321876e5;
			s_box3[118]<= 32'h96e7365c;
			s_box3[119]<= 32'h96b52815;
			s_box3[120]<= 32'h02919d67;
			s_box3[121]<= 32'h6f62b721;
			s_box3[122]<= 32'h322f9862;
			s_box3[123]<= 32'h9407760d;
			s_box3[124]<= 32'h875f12a2;
			s_box3[125]<= 32'h9674994d;
			s_box3[126]<= 32'h27f311c1;
			s_box3[127]<= 32'h445171af;
			s_box3[128]<= 32'h0d09222c;
			s_box3[129]<= 32'h986427b3;
			s_box3[130]<= 32'h68962b8c;
			s_box3[131]<= 32'h9f168f51;
			s_box3[132]<= 32'h8ba8122c;
			s_box3[133]<= 32'h15f33668;
			s_box3[134]<= 32'h6109439f;
			s_box3[135]<= 32'h991c4c16;
			s_box3[136]<= 32'h07d9f783;
			s_box3[137]<= 32'h9c762744;
			s_box3[138]<= 32'h79949d1c;
			s_box3[139]<= 32'h017596a7;
			s_box3[140]<= 32'h74c803d9;
			s_box3[141]<= 32'h2565615f;
			s_box3[142]<= 32'h1d670606;
			s_box3[143]<= 32'h69655928;
			s_box3[144]<= 32'h70a8276f;
			s_box3[145]<= 32'h5c246f91;
			s_box3[146]<= 32'h5f69a528;
			s_box3[147]<= 32'h8674995b;
			s_box3[148]<= 32'h80d5d71c;
			s_box3[149]<= 32'h5c197992;
			s_box3[150]<= 32'h567922d3;
			s_box3[151]<= 32'h5c3327d1;
			s_box3[152]<= 32'h40c952c7;
			s_box3[153]<= 32'h52a67744;
			s_box3[154]<= 32'h6a908906;
			s_box3[155]<= 32'h42636952;
			s_box3[156]<= 32'h508a65b7;
			s_box3[157]<= 32'h2499d7a2;
			s_box3[158]<= 32'h7d922572;
			s_box3[159]<= 32'h0491953f;
			s_box3[160]<= 32'h52495c61;
			s_box3[161]<= 32'h40c88599;
			s_box3[162]<= 32'h7207aef0;
			s_box3[163]<= 32'h98d169d5;
			s_box3[164]<= 32'h45455a73;
			s_box3[165]<= 32'h9658257a;
			s_box3[166]<= 32'h089c8915;
			s_box3[167]<= 32'h4223b24f;
			s_box3[168]<= 32'h98c7e39a;
			s_box3[169]<= 32'h2b96312a;
			s_box3[170]<= 32'h75b63e79;
			s_box3[171]<= 32'h58bfb5a0;
			s_box3[172]<= 32'h9750c3a9;
			s_box3[173]<= 32'h22c8c459;
			s_box3[174]<= 32'h76b32549;
			s_box3[175]<= 32'h8cdc3a36;
			s_box3[176]<= 32'h89151608;
			s_box3[177]<= 32'h2f87c582;
			s_box3[178]<= 32'h196291b1;
			s_box3[179]<= 32'h5b056ef8;
			s_box3[180]<= 32'h9c7a08b5;
			s_box3[181]<= 32'h84c8515f;
			s_box3[182]<= 32'h0d62b95b;
			s_box3[183]<= 32'h662a0c71;
			s_box3[184]<= 32'h56722237;
			s_box3[185]<= 32'h6f5f849c;
			s_box3[186]<= 32'h262a3641;
			s_box3[187]<= 32'h4b34b631;
			s_box3[188]<= 32'h4f923c72;
			s_box3[189]<= 32'h4f989c1c;
			s_box3[190]<= 32'h5c6b4594;
			s_box3[191]<= 32'h27f29910;
			s_box3[192]<= 32'h21571217;
			s_box3[193]<= 32'h45455a73;
			s_box3[194]<= 32'h804d9561;
			s_box3[195]<= 32'h515792c8;
			s_box3[196]<= 32'h567922d3;
			s_box3[197]<= 32'h706b4765;
			s_box3[198]<= 32'h5a2971d5;
			s_box3[199]<= 32'h5f74f74d;
			s_box3[200]<= 32'h82728952;
			s_box3[201]<= 32'h217c2a71;
			s_box3[202]<= 32'h321876e5;
			s_box3[203]<= 32'h96e7365c;
			s_box3[204]<= 32'h96b52815;
			s_box3[205]<= 32'h02919d67;
			s_box3[206]<= 32'h6f62b721;
			s_box3[207]<= 32'h322f9862;
			s_box3[208]<= 32'h9407760d;
			s_box3[209]<= 32'h875f12a2;
			s_box3[210]<= 32'h9674994d;
			s_box3[211]<= 32'h27f311c1;
			s_box3[212]<= 32'h445171af;
			s_box3[213]<= 32'h0d09222c;
			s_box3[214]<= 32'h986427b3;
			s_box3[215]<= 32'h68962b8c;
			s_box3[216]<= 32'h9f168f51;
			s_box3[217]<= 32'h8ba8122c;
			s_box3[218]<= 32'h15f33668;
			s_box3[219]<= 32'h6109439f;
			s_box3[220]<= 32'h991c4c16;
			s_box3[221]<= 32'h07d9f783;
			s_box3[222]<= 32'h9c762744;
			s_box3[223]<= 32'h79949d1c;
			s_box3[224]<= 32'h017596a7;
			s_box3[225]<= 32'h74c803d9;
			s_box3[226]<= 32'h2565615f;
			s_box3[227]<= 32'h1d670606;
			s_box3[228]<= 32'h69655928;
			s_box3[229]<= 32'h70a8276f;
			s_box3[230]<= 32'h5c246f91;
			s_box3[231]<= 32'h5f69a528;
			s_box3[232]<= 32'h8674995b;
			s_box3[233]<= 32'h80d5d71c;
			s_box3[234]<= 32'h5c197992;
			s_box3[235]<= 32'h567922d3;
			s_box3[236]<= 32'h5c3327d1;
			s_box3[237]<= 32'h40c952c7;
			s_box3[238]<= 32'h52a67744;
			s_box3[239]<= 32'h6a908906;
			s_box3[240]<= 32'h42636952;
			s_box3[241]<= 32'h508a65b7;
			s_box3[242]<= 32'h2499d7a2;
			s_box3[243]<= 32'h7d922572;
			s_box3[244]<= 32'h0491953f;
			s_box3[245]<= 32'h52495c61;
			s_box3[246]<= 32'h40c88599;
			s_box3[247]<= 32'h7207aef0;
			s_box3[248]<= 32'h98d169d5;
			s_box3[249]<= 32'h45455a73;
			s_box3[250]<= 32'h9658257a;
			s_box3[251]<= 32'h089c8915;
			s_box3[252]<= 32'h4223b24f;
			s_box3[253]<= 32'h98c7e39a;
			s_box3[254]<= 32'h2b96312a;
			s_box3[255]<= 32'h75b63e79;

            right <= 0;
            left  <= 0;
            temp  <= 0;

            round <= 0;

            DECRYPT_DONE  <= 0;
            decryptedtext <= 64'h0;

            state <= IDLE;

        end else begin
            case (state)

                IDLE: begin
                    if (!start)
                        state <= INIT;
                    else
                        state <= TRANSITION;
                end

                TRANSITION: begin
                    if (start && !DECRYPT_DONE) begin
                        left  <= ciphertext[63:32];
                        right <= ciphertext[31:0];
                        round <= 15;
                        state <= ENCRYPT_UNDO;
                    end else begin
                        state <= IDLE;
                    end
                end

                INIT: begin
                    init  <= 1;
                    state <= IDLE;
                end

                ENCRYPT_UNDO: begin
                    left  <= ciphertext[63:32] ^ p_array[16];
                    right <= ciphertext[31:0]  ^ p_array[17];
                    state <= DECRYPT_RIGHT;
                end

                DECRYPT_RIGHT: begin
                    temp  <= right;
                    right <= left ^ p_array[round];
                    state <= DECRYPT_LEFT;
                end

                DECRYPT_LEFT: begin
                    left  <= temp ^ F(left);
                    round <= round - 1;

                    if (round == 0)
                        state <= DONE;
                    else
                        state <= DECRYPT_RIGHT;
                end

                DONE: begin
                    decryptedtext <= {right, left};
                    DECRYPT_DONE  <= 1;
                    state         <= IDLE;
                end

                default: state <= IDLE;

            endcase
        end
    end

endmodule
